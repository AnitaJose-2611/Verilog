module NOTGate(
  input a,
  output out
);
  assign out = ~a;
endmodule
